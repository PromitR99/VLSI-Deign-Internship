module full_subtractor_tb();

  reg   a,b,bin;
  wire  diff,borrow;
 
  integer i;

  //Instantiate the full adder
  full_subtractor DUT(.a(a), .b(b), .b_in(bin), .diff(diff), .borrow(borrow));

  initial 
  begin
    a   = 1'b0;
    b   = 1'b0;
    bin = 1'b0;
  end

  initial
  begin 
    for (i=0;i<8;i=i+1)
    begin
      {a,b,bin}=i;
      #10;
    end
  end

  initial $monitor("Input a=%b, b=%b, c=%b, Output sum =%b, carry=%b",
                  a,b,bin,diff,borrow);

  initial #100 $finish;

endmodule